//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat May 24 14:04:13 2025
//-------------------------------------------
// ----- Verilog module for fpga_top -----
module fpga_top(prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:11] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:8] cbx_1__0__0_chanx_left_out;
wire [0:8] cbx_1__0__0_chanx_right_out;
wire [0:8] cbx_1__0__1_chanx_left_out;
wire [0:8] cbx_1__0__1_chanx_right_out;
wire [0:8] cbx_1__0__2_chanx_left_out;
wire [0:8] cbx_1__0__2_chanx_right_out;
wire [0:8] cbx_1__1__0_chanx_left_out;
wire [0:8] cbx_1__1__0_chanx_right_out;
wire [0:8] cbx_1__1__1_chanx_left_out;
wire [0:8] cbx_1__1__1_chanx_right_out;
wire [0:8] cbx_1__1__2_chanx_left_out;
wire [0:8] cbx_1__1__2_chanx_right_out;
wire [0:8] cbx_1__1__3_chanx_left_out;
wire [0:8] cbx_1__1__3_chanx_right_out;
wire [0:8] cbx_1__1__4_chanx_left_out;
wire [0:8] cbx_1__1__4_chanx_right_out;
wire [0:8] cbx_1__1__5_chanx_left_out;
wire [0:8] cbx_1__1__5_chanx_right_out;
wire [0:8] cbx_1__3__0_chanx_left_out;
wire [0:8] cbx_1__3__0_chanx_right_out;
wire [0:8] cbx_1__3__1_chanx_left_out;
wire [0:8] cbx_1__3__1_chanx_right_out;
wire [0:8] cbx_1__3__2_chanx_left_out;
wire [0:8] cbx_1__3__2_chanx_right_out;
wire [0:8] cby_0__1__0_chany_bottom_out;
wire [0:8] cby_0__1__0_chany_top_out;
wire [0:8] cby_0__1__1_chany_bottom_out;
wire [0:8] cby_0__1__1_chany_top_out;
wire [0:8] cby_0__1__2_chany_bottom_out;
wire [0:8] cby_0__1__2_chany_top_out;
wire [0:8] cby_1__1__0_chany_bottom_out;
wire [0:8] cby_1__1__0_chany_top_out;
wire [0:8] cby_1__1__1_chany_bottom_out;
wire [0:8] cby_1__1__1_chany_top_out;
wire [0:8] cby_1__1__2_chany_bottom_out;
wire [0:8] cby_1__1__2_chany_top_out;
wire [0:8] cby_1__1__3_chany_bottom_out;
wire [0:8] cby_1__1__3_chany_top_out;
wire [0:8] cby_1__1__4_chany_bottom_out;
wire [0:8] cby_1__1__4_chany_top_out;
wire [0:8] cby_1__1__5_chany_bottom_out;
wire [0:8] cby_1__1__5_chany_top_out;
wire [0:8] cby_3__1__0_chany_bottom_out;
wire [0:8] cby_3__1__0_chany_top_out;
wire [0:8] cby_3__1__1_chany_bottom_out;
wire [0:8] cby_3__1__1_chany_top_out;
wire [0:8] cby_3__1__2_chany_bottom_out;
wire [0:8] cby_3__1__2_chany_top_out;
wire [0:8] sb_0__0__0_chanx_right_out;
wire [0:8] sb_0__0__0_chany_top_out;
wire [0:8] sb_0__1__0_chanx_right_out;
wire [0:8] sb_0__1__0_chany_bottom_out;
wire [0:8] sb_0__1__0_chany_top_out;
wire [0:8] sb_0__1__1_chanx_right_out;
wire [0:8] sb_0__1__1_chany_bottom_out;
wire [0:8] sb_0__1__1_chany_top_out;
wire [0:8] sb_0__3__0_chanx_right_out;
wire [0:8] sb_0__3__0_chany_bottom_out;
wire [0:8] sb_1__0__0_chanx_left_out;
wire [0:8] sb_1__0__0_chanx_right_out;
wire [0:8] sb_1__0__0_chany_top_out;
wire [0:8] sb_1__0__1_chanx_left_out;
wire [0:8] sb_1__0__1_chanx_right_out;
wire [0:8] sb_1__0__1_chany_top_out;
wire [0:8] sb_1__1__0_chanx_left_out;
wire [0:8] sb_1__1__0_chanx_right_out;
wire [0:8] sb_1__1__0_chany_bottom_out;
wire [0:8] sb_1__1__0_chany_top_out;
wire [0:8] sb_1__1__1_chanx_left_out;
wire [0:8] sb_1__1__1_chanx_right_out;
wire [0:8] sb_1__1__1_chany_bottom_out;
wire [0:8] sb_1__1__1_chany_top_out;
wire [0:8] sb_1__1__2_chanx_left_out;
wire [0:8] sb_1__1__2_chanx_right_out;
wire [0:8] sb_1__1__2_chany_bottom_out;
wire [0:8] sb_1__1__2_chany_top_out;
wire [0:8] sb_1__1__3_chanx_left_out;
wire [0:8] sb_1__1__3_chanx_right_out;
wire [0:8] sb_1__1__3_chany_bottom_out;
wire [0:8] sb_1__1__3_chany_top_out;
wire [0:8] sb_1__3__0_chanx_left_out;
wire [0:8] sb_1__3__0_chanx_right_out;
wire [0:8] sb_1__3__0_chany_bottom_out;
wire [0:8] sb_1__3__1_chanx_left_out;
wire [0:8] sb_1__3__1_chanx_right_out;
wire [0:8] sb_1__3__1_chany_bottom_out;
wire [0:8] sb_3__0__0_chanx_left_out;
wire [0:8] sb_3__0__0_chany_top_out;
wire [0:8] sb_3__1__0_chanx_left_out;
wire [0:8] sb_3__1__0_chany_bottom_out;
wire [0:8] sb_3__1__0_chany_top_out;
wire [0:8] sb_3__1__1_chanx_left_out;
wire [0:8] sb_3__1__1_chany_bottom_out;
wire [0:8] sb_3__1__1_chany_top_out;
wire [0:8] sb_3__3__0_chanx_left_out;
wire [0:8] sb_3__3__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__3__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[1]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__3__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[2]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__3__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_right grid_io_right_4__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[3]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_4__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[4]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_4__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[5]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[6]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[7]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[9]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[10]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[11]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_3__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_3__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_3__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(ccff_tail));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:8]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:8]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(sb_0__3__0_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__3_ sb_0__3_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__3__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__3__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__3__0_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__3__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_2__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__3_ sb_1__3_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__3__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__3__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__3__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__3__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__3__0_ccff_tail));

	sb_1__3_ sb_2__3_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__3__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__3__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__3__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__3__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__3__1_ccff_tail));

	sb_3__0_ sb_3__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_3__0__0_chany_top_out[0:8]),
		.chanx_left_out(sb_3__0__0_chanx_left_out[0:8]),
		.ccff_tail(sb_3__0__0_ccff_tail));

	sb_3__1_ sb_3__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_3__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_3__1__0_chany_top_out[0:8]),
		.chany_bottom_out(sb_3__1__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_3__1__0_chanx_left_out[0:8]),
		.ccff_tail(sb_3__1__0_ccff_tail));

	sb_3__1_ sb_3__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_3__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_3__1__1_chany_top_out[0:8]),
		.chany_bottom_out(sb_3__1__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_3__1__1_chanx_left_out[0:8]),
		.ccff_tail(sb_3__1__1_ccff_tail));

	sb_3__3_ sb_3__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_3__3__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_3__3__0_chanx_left_out[0:8]),
		.ccff_tail(sb_3__3__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_3__0__0_chanx_left_out[0:8]),
		.ccff_head(sb_3__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_2__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:8]),
		.chanx_right_in(sb_3__1__0_chanx_left_out[0:8]),
		.ccff_head(sb_3__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:8]),
		.chanx_right_in(sb_3__1__1_chanx_left_out[0:8]),
		.ccff_head(sb_3__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__3_ cbx_1__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__3__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__3__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__0_ccff_tail));

	cbx_1__3_ cbx_2__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__3__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__3__1_ccff_tail),
		.chanx_left_out(cbx_1__3__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__3__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__1_ccff_tail));

	cbx_1__3_ cbx_3__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_3__3__0_chanx_left_out[0:8]),
		.ccff_head(sb_3__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__3__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__2_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:8]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_0__3__0_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_1__3__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:8]),
		.chany_top_in(sb_1__3__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_3__1_ cby_3__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_3__1__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_3__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_3__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_3__1__0_ccff_tail));

	cby_3__1_ cby_3__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_3__1__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_bottom_out(cby_3__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_3__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_3__1__1_ccff_tail));

	cby_3__1_ cby_3__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_3__3__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_3__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_3__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_3__1__2_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----




